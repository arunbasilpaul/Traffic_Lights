library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package TRAFFIC_TYPES is
	type TRAFFIC_LIGHT is (RED, GREEN, YELLOW, PENDING);
end package TRAFFIC_TYPES; 